module main

import dbops

fn main() {
	dbops.connect_db()
}